module layer1_tcbcnn_121_25x64x10
(
    input clk,
    input rst,
    input [1728-1:0] layer_in,
    input valid,
    output  reg ready,
    output [36*10-1:0] layer_out
);
parameter DATA_WIDTH = 36;
parameter INPUT_DATA_CNT   =   64;
reg    signed [27-1:0]  in_buffer[0:INPUT_DATA_CNT-1];
genvar j;
generate
for(j=0;j<INPUT_DATA_CNT;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=layer_in[j*27+26:j*27+0];
                    end
            end
    end
endgenerate
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight0;
assign in_buffer_weight0=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<4))-(0+(in_buffer[2]<<0)+(in_buffer[2]<<2)+(in_buffer[2]<<4)+(in_buffer[2]<<5))+(0+(in_buffer[3]<<0)+(in_buffer[3]<<2)+(in_buffer[3]<<4)+(in_buffer[3]<<6))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2))+(0+(in_buffer[5]<<0)+(in_buffer[5]<<1))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<4)+(in_buffer[6]<<6))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<4)+(in_buffer[7]<<5))+(0+(in_buffer[8]<<0)+(in_buffer[8]<<3)+(in_buffer[8]<<5))-(0-(in_buffer[9]<<3)+(in_buffer[9]<<6))+(0-(in_buffer[10]<<1)+(in_buffer[10]<<6))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<2)+(in_buffer[11]<<3))+(0+(in_buffer[12]<<3)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<1)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<3))+(0-(in_buffer[15]<<1)+(in_buffer[15]<<4))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<3)+(in_buffer[16]<<5)+(in_buffer[16]<<6))-(0+(in_buffer[17]<<4)+(in_buffer[17]<<7))+(0+(in_buffer[18]<<0)+(in_buffer[18]<<5))+(0-(in_buffer[19]<<1)-(in_buffer[19]<<3)+(in_buffer[19]<<6))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<3)+(in_buffer[21]<<4))-(0-(in_buffer[22]<<0)+(in_buffer[22]<<3))-(0+(in_buffer[23]<<4)+(in_buffer[23]<<5))+(0-(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<4))-(0-(in_buffer[25]<<3)+(in_buffer[25]<<5)+(in_buffer[25]<<6))-(0+(in_buffer[26]<<0)+(in_buffer[26]<<2)-(in_buffer[26]<<4)+(in_buffer[26]<<7))+(0-(in_buffer[27]<<2)+(in_buffer[27]<<5))+(0-(in_buffer[28]<<0)-(in_buffer[28]<<3)+(in_buffer[28]<<6)+(in_buffer[28]<<7))-(0+(in_buffer[29]<<0)+(in_buffer[29]<<2)-(in_buffer[29]<<4)+(in_buffer[29]<<7))-(0+(in_buffer[30]<<0)+(in_buffer[30]<<2)+(in_buffer[30]<<5))+(0+(in_buffer[31]<<2)+(in_buffer[31]<<3))+(0+(in_buffer[32]<<0)+(in_buffer[32]<<2)+(in_buffer[32]<<4))+(0+(in_buffer[33]<<6))+(0+(in_buffer[34]<<0)+(in_buffer[34]<<3))-(0+(in_buffer[35]<<2)+(in_buffer[35]<<4)+(in_buffer[35]<<6))-(0+(in_buffer[36]<<1)+(in_buffer[36]<<3)+(in_buffer[36]<<6)+(in_buffer[36]<<7))-(0-(in_buffer[37]<<0)+(in_buffer[37]<<4))-(0-(in_buffer[38]<<0)+(in_buffer[38]<<7))-(0-(in_buffer[39]<<2)-(in_buffer[39]<<4)+(in_buffer[39]<<7))-(0+(in_buffer[40]<<0)+(in_buffer[40]<<2))+(0+(in_buffer[41]<<0)+(in_buffer[41]<<1)+(in_buffer[41]<<4)+(in_buffer[41]<<5))+(0+(in_buffer[42]<<0)+(in_buffer[42]<<5))-(0+(in_buffer[43]<<1)+(in_buffer[43]<<2))+(0+(in_buffer[44]<<0)+(in_buffer[44]<<2))-(0-(in_buffer[45]<<2)+(in_buffer[45]<<8))+(0+(in_buffer[46]<<0)+(in_buffer[46]<<1)+(in_buffer[46]<<6))-(0+(in_buffer[47]<<1))+(0+(in_buffer[48]<<0))-(0-(in_buffer[49]<<1)+(in_buffer[49]<<4)+(in_buffer[49]<<5))-(0-(in_buffer[50]<<1)-(in_buffer[50]<<4)+(in_buffer[50]<<6)+(in_buffer[50]<<7))-(0+(in_buffer[51]<<0)+(in_buffer[51]<<1)+(in_buffer[51]<<5))+(0+(in_buffer[52]<<0)+(in_buffer[52]<<1)+(in_buffer[52]<<7))+(0-(in_buffer[53]<<1)+(in_buffer[53]<<4)+(in_buffer[53]<<6))-(0+(in_buffer[54]<<3)+(in_buffer[54]<<6))+(0-(in_buffer[55]<<0)+(in_buffer[55]<<2)+(in_buffer[55]<<3)+(in_buffer[55]<<6))+(0+(in_buffer[56]<<4)+(in_buffer[56]<<6))-(0+(in_buffer[57]<<0)+(in_buffer[57]<<3)+(in_buffer[57]<<5))+(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)+(in_buffer[58]<<3))-(0-(in_buffer[59]<<0)+(in_buffer[59]<<2)+(in_buffer[59]<<3))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)+(in_buffer[60]<<5)+(in_buffer[60]<<6))-(0+(in_buffer[61]<<0)+(in_buffer[61]<<3))-(0-(in_buffer[62]<<1)-(in_buffer[62]<<3)+(in_buffer[62]<<6))+(0+(in_buffer[63]<<4)+(in_buffer[63]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight1;
assign in_buffer_weight1=0+(0+(in_buffer[0]<<4))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<1))+(0+(in_buffer[2]<<1)+(in_buffer[2]<<2))-(0+(in_buffer[3]<<2)+(in_buffer[3]<<6))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<6))+(0+(in_buffer[5]<<0)+(in_buffer[5]<<2)+(in_buffer[5]<<3))-(0-(in_buffer[6]<<1)+(in_buffer[6]<<4))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<2))-(0+(in_buffer[8]<<0)+(in_buffer[8]<<1)+(in_buffer[8]<<5)+(in_buffer[8]<<6))+(0+(in_buffer[9]<<0)-(in_buffer[9]<<2)+(in_buffer[9]<<6))-(0-(in_buffer[10]<<0)+(in_buffer[10]<<4)+(in_buffer[10]<<6))+(0+(in_buffer[11]<<0)+(in_buffer[11]<<1)+(in_buffer[11]<<4)+(in_buffer[11]<<7))+(0+(in_buffer[12]<<2)+(in_buffer[12]<<5)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<1)+(in_buffer[13]<<3)+(in_buffer[13]<<5))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3))+(0+(in_buffer[16]<<0)-(in_buffer[16]<<2)+(in_buffer[16]<<4)+(in_buffer[16]<<5))+(0+(in_buffer[17]<<4)+(in_buffer[17]<<5))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<2)+(in_buffer[19]<<3))-(0+(in_buffer[20]<<0)+(in_buffer[20]<<5)+(in_buffer[20]<<6))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<2)+(in_buffer[21]<<5)+(in_buffer[21]<<6))+(0-(in_buffer[22]<<1)+(in_buffer[22]<<5))-(0-(in_buffer[23]<<0)-(in_buffer[23]<<3)+(in_buffer[23]<<5)+(in_buffer[23]<<6))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<6))+(0-(in_buffer[25]<<0)+(in_buffer[25]<<2)+(in_buffer[25]<<3))+(0+(in_buffer[26]<<1)+(in_buffer[26]<<3)+(in_buffer[26]<<5))-(0+(in_buffer[27]<<1)+(in_buffer[27]<<3)+(in_buffer[27]<<5)+(in_buffer[27]<<6))+(0+(in_buffer[28]<<3))-(0-(in_buffer[29]<<0)+(in_buffer[29]<<3))-(0-(in_buffer[31]<<0)+(in_buffer[31]<<3))+(0-(in_buffer[32]<<0)-(in_buffer[32]<<2)+(in_buffer[32]<<5))+(0+(in_buffer[33]<<0)+(in_buffer[33]<<2)+(in_buffer[33]<<4)+(in_buffer[33]<<5))-(0+(in_buffer[34]<<0)+(in_buffer[34]<<5)+(in_buffer[34]<<6))-(0+(in_buffer[35]<<0)+(in_buffer[35]<<3))+(0+(in_buffer[36]<<0)+(in_buffer[36]<<1))-(0+(in_buffer[37]<<0)+(in_buffer[37]<<1)+(in_buffer[37]<<6))+(0+(in_buffer[38]<<0))-(0-(in_buffer[39]<<0)+(in_buffer[39]<<4)+(in_buffer[39]<<5))-(0+(in_buffer[40]<<2)+(in_buffer[40]<<3))+(0+(in_buffer[41]<<1)+(in_buffer[41]<<3)+(in_buffer[41]<<5)+(in_buffer[41]<<6))+(0+(in_buffer[42]<<0)+(in_buffer[42]<<2)+(in_buffer[42]<<4)+(in_buffer[42]<<5))+(0+(in_buffer[43]<<2)-(in_buffer[43]<<4)+(in_buffer[43]<<7))-(0-(in_buffer[44]<<1)+(in_buffer[44]<<4)+(in_buffer[44]<<6)+(in_buffer[44]<<7))+(0+(in_buffer[45]<<0)+(in_buffer[45]<<2)+(in_buffer[45]<<5)+(in_buffer[45]<<6))+(0+(in_buffer[46]<<0)+(in_buffer[46]<<2)+(in_buffer[46]<<5)+(in_buffer[46]<<6))-(0+(in_buffer[47]<<0))-(0-(in_buffer[48]<<0)-(in_buffer[48]<<3)+(in_buffer[48]<<5)+(in_buffer[48]<<6))-(0+(in_buffer[49]<<0)+(in_buffer[49]<<2)+(in_buffer[49]<<4)+(in_buffer[49]<<6))+(0+(in_buffer[50]<<1)+(in_buffer[50]<<3)+(in_buffer[50]<<6))+(0+(in_buffer[51]<<1)+(in_buffer[51]<<2)+(in_buffer[51]<<5))-(0+(in_buffer[52]<<2)+(in_buffer[52]<<3)+(in_buffer[52]<<6))-(0-(in_buffer[53]<<1)+(in_buffer[53]<<4)+(in_buffer[53]<<5))+(0+(in_buffer[54]<<4)+(in_buffer[54]<<5))-(0-(in_buffer[55]<<4)+(in_buffer[55]<<7))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<1)-(in_buffer[56]<<4)+(in_buffer[56]<<6)+(in_buffer[56]<<7))+(0+(in_buffer[57]<<1)+(in_buffer[57]<<3))+(0+(in_buffer[58]<<2)+(in_buffer[58]<<5))+(0+(in_buffer[59]<<0)+(in_buffer[59]<<1))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)+(in_buffer[60]<<4))+(0+(in_buffer[61]<<0)+(in_buffer[61]<<4)+(in_buffer[61]<<6))+(0-(in_buffer[62]<<0)-(in_buffer[62]<<3)+(in_buffer[62]<<7))-(0+(in_buffer[63]<<1)+(in_buffer[63]<<3)+(in_buffer[63]<<5)+(in_buffer[63]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight2;
assign in_buffer_weight2=0+(0-(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3))+(0-(in_buffer[1]<<2)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<2)+(in_buffer[2]<<4))-(0+(in_buffer[3]<<1))+(0+(in_buffer[4]<<1)-(in_buffer[4]<<3)+(in_buffer[4]<<6))+(0+(in_buffer[5]<<2)+(in_buffer[5]<<3))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<1)+(in_buffer[6]<<6))+(0+(in_buffer[7]<<2)+(in_buffer[7]<<4))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<8))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<3))-(0-(in_buffer[10]<<0)+(in_buffer[10]<<6))+(0+(in_buffer[11]<<0)-(in_buffer[11]<<2)+(in_buffer[11]<<5))+(0+(in_buffer[12]<<1)-(in_buffer[12]<<3)+(in_buffer[12]<<6))+(0+(in_buffer[13]<<4))+(0+(in_buffer[14]<<0)+(in_buffer[14]<<2)+(in_buffer[14]<<3))-(0+(in_buffer[15]<<3))-(0+(in_buffer[16]<<0)+(in_buffer[16]<<3)+(in_buffer[16]<<5))+(0-(in_buffer[17]<<1)+(in_buffer[17]<<6))+(0+(in_buffer[18]<<1)-(in_buffer[18]<<3)+(in_buffer[18]<<6))+(0-(in_buffer[19]<<0)-(in_buffer[19]<<4)+(in_buffer[19]<<7))-(0+(in_buffer[20]<<0)-(in_buffer[20]<<3)+(in_buffer[20]<<6))-(0+(in_buffer[21]<<2)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<3)+(in_buffer[22]<<5))-(0+(in_buffer[23]<<0)-(in_buffer[23]<<2)+(in_buffer[23]<<5)+(in_buffer[23]<<6))-(0+(in_buffer[24]<<0)+(in_buffer[24]<<2))+(0+(in_buffer[25]<<0)+(in_buffer[25]<<2)+(in_buffer[25]<<4)+(in_buffer[25]<<5))-(0+(in_buffer[26]<<0)-(in_buffer[26]<<2)+(in_buffer[26]<<4)+(in_buffer[26]<<5))+(0+(in_buffer[27]<<3))+(0-(in_buffer[28]<<0)+(in_buffer[28]<<3)+(in_buffer[28]<<5))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<2)+(in_buffer[29]<<3))-(0+(in_buffer[30]<<3)+(in_buffer[30]<<4)+(in_buffer[30]<<7))-(0+(in_buffer[31]<<3))-(0+(in_buffer[32]<<1)+(in_buffer[32]<<5))-(0+(in_buffer[33]<<0)-(in_buffer[33]<<3)+(in_buffer[33]<<5)+(in_buffer[33]<<6))-(0-(in_buffer[34]<<0)-(in_buffer[34]<<3)+(in_buffer[34]<<6))-(0-(in_buffer[35]<<0)-(in_buffer[35]<<2)+(in_buffer[35]<<5)+(in_buffer[35]<<7))+(0-(in_buffer[36]<<1)+(in_buffer[36]<<4)+(in_buffer[36]<<5))-(0-(in_buffer[37]<<0)-(in_buffer[37]<<2)-(in_buffer[37]<<4)+(in_buffer[37]<<7))+(0+(in_buffer[38]<<0)+(in_buffer[38]<<3)+(in_buffer[38]<<4)+(in_buffer[38]<<7))-(0+(in_buffer[39]<<2)+(in_buffer[39]<<3)+(in_buffer[39]<<6)+(in_buffer[39]<<7))-(0+(in_buffer[40]<<1)+(in_buffer[40]<<3))-(0+(in_buffer[41]<<5))-(0+(in_buffer[42]<<3))-(0+(in_buffer[43]<<2)+(in_buffer[43]<<4))-(0+(in_buffer[44]<<0)+(in_buffer[44]<<3)+(in_buffer[44]<<4))+(0+(in_buffer[45]<<0)+(in_buffer[45]<<3)+(in_buffer[45]<<5))+(0+(in_buffer[46]<<1)+(in_buffer[46]<<4))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<3))-(0-(in_buffer[48]<<1)-(in_buffer[48]<<3)+(in_buffer[48]<<6)+(in_buffer[48]<<7))-(0+(in_buffer[49]<<2))+(0+(in_buffer[50]<<1)+(in_buffer[50]<<2))+(0-(in_buffer[51]<<0)+(in_buffer[51]<<4)+(in_buffer[51]<<5))+(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<5)+(in_buffer[52]<<6))+(0-(in_buffer[53]<<0)+(in_buffer[53]<<4)+(in_buffer[53]<<5))+(0-(in_buffer[54]<<0)+(in_buffer[54]<<4)+(in_buffer[54]<<5))+(0-(in_buffer[55]<<0)+(in_buffer[55]<<2)+(in_buffer[55]<<3))+(0+(in_buffer[56]<<0)+(in_buffer[56]<<4))-(0+(in_buffer[57]<<1)+(in_buffer[57]<<2))+(0-(in_buffer[58]<<1)+(in_buffer[58]<<4)+(in_buffer[58]<<6))+(0+(in_buffer[59]<<2))+(0+(in_buffer[60]<<2))-(0+(in_buffer[61]<<2)+(in_buffer[61]<<4)+(in_buffer[61]<<6))+(0+(in_buffer[62]<<0)+(in_buffer[62]<<1))-(0-(in_buffer[63]<<2)+(in_buffer[63]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight3;
assign in_buffer_weight3=0+(0+(in_buffer[0]<<2)+(in_buffer[0]<<3))-(0+(in_buffer[1]<<4)+(in_buffer[1]<<6))+(0-(in_buffer[2]<<0)+(in_buffer[2]<<2)+(in_buffer[2]<<3))+(0+(in_buffer[3]<<2)+(in_buffer[3]<<3))+(0+(in_buffer[4]<<0)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<1)+(in_buffer[5]<<4))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<3)+(in_buffer[6]<<5))-(0+(in_buffer[7]<<4))+(0+(in_buffer[8]<<1)+(in_buffer[8]<<2)+(in_buffer[8]<<5))-(0+(in_buffer[9]<<0)-(in_buffer[9]<<3)+(in_buffer[9]<<6))-(0+(in_buffer[10]<<1)+(in_buffer[10]<<4))-(0-(in_buffer[11]<<0)+(in_buffer[11]<<3))-(0+(in_buffer[12]<<2)+(in_buffer[12]<<6))+(0+(in_buffer[13]<<0)+(in_buffer[13]<<3))-(0+(in_buffer[14]<<0)+(in_buffer[14]<<2))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3))+(0+(in_buffer[16]<<2)+(in_buffer[16]<<4)+(in_buffer[16]<<5))-(0-(in_buffer[17]<<0)+(in_buffer[17]<<2)+(in_buffer[17]<<3)+(in_buffer[17]<<6))-(0+(in_buffer[18]<<3)+(in_buffer[18]<<4))-(0-(in_buffer[19]<<0)-(in_buffer[19]<<4)+(in_buffer[19]<<7))+(0+(in_buffer[20]<<2)+(in_buffer[20]<<4))-(0+(in_buffer[21]<<0)-(in_buffer[21]<<2)+(in_buffer[21]<<5))+(0+(in_buffer[22]<<3)+(in_buffer[22]<<5))+(0-(in_buffer[23]<<2)+(in_buffer[23]<<6))+(0-(in_buffer[24]<<1)+(in_buffer[24]<<3)+(in_buffer[24]<<4))+(0+(in_buffer[25]<<0)+(in_buffer[25]<<6))+(0+(in_buffer[26]<<1))-(0-(in_buffer[27]<<0)+(in_buffer[27]<<3)+(in_buffer[27]<<5))-(0+(in_buffer[28]<<3)+(in_buffer[28]<<5))-(0-(in_buffer[29]<<0)+(in_buffer[29]<<7))+(0+(in_buffer[30]<<1)+(in_buffer[30]<<3)+(in_buffer[30]<<4))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<2)+(in_buffer[31]<<3))-(0+(in_buffer[32]<<0)+(in_buffer[32]<<2)+(in_buffer[32]<<4))-(0-(in_buffer[33]<<2)-(in_buffer[33]<<4)+(in_buffer[33]<<6)+(in_buffer[33]<<7))+(0+(in_buffer[34]<<1)+(in_buffer[34]<<5))-(0-(in_buffer[35]<<1)+(in_buffer[35]<<5))+(0+(in_buffer[36]<<1)+(in_buffer[36]<<3)+(in_buffer[36]<<4))-(0+(in_buffer[37]<<0)+(in_buffer[37]<<1)+(in_buffer[37]<<6))+(0+(in_buffer[39]<<5)+(in_buffer[39]<<6))+(0+(in_buffer[40]<<2))-(0+(in_buffer[41]<<2)+(in_buffer[41]<<6))+(0-(in_buffer[42]<<0)+(in_buffer[42]<<2)+(in_buffer[42]<<3))+(0-(in_buffer[43]<<0)+(in_buffer[43]<<4))+(0+(in_buffer[44]<<0))+(0+(in_buffer[45]<<2)+(in_buffer[45]<<5))+(0-(in_buffer[46]<<1)+(in_buffer[46]<<4))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<1))+(0-(in_buffer[48]<<0)+(in_buffer[48]<<2)+(in_buffer[48]<<3))+(0+(in_buffer[50]<<0)+(in_buffer[50]<<1)+(in_buffer[50]<<5))+(0-(in_buffer[51]<<1)+(in_buffer[51]<<5))-(0+(in_buffer[52]<<0)+(in_buffer[52]<<4))+(0+(in_buffer[53]<<0)+(in_buffer[53]<<6))-(0+(in_buffer[54]<<3)+(in_buffer[54]<<5))+(0+(in_buffer[55]<<1)+(in_buffer[55]<<5))+(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<3))-(0-(in_buffer[57]<<1)+(in_buffer[57]<<5))+(0-(in_buffer[58]<<2)+(in_buffer[58]<<4)+(in_buffer[58]<<5))-(0+(in_buffer[59]<<3))+(0+(in_buffer[60]<<0)+(in_buffer[60]<<1)+(in_buffer[60]<<5))+(0+(in_buffer[61]<<4))-(0+(in_buffer[62]<<5)+(in_buffer[62]<<6))+(0-(in_buffer[63]<<0)+(in_buffer[63]<<3)+(in_buffer[63]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight4;
assign in_buffer_weight4=0+(0+(in_buffer[0]<<2))+(0+(in_buffer[1]<<0)-(in_buffer[1]<<3)+(in_buffer[1]<<6))+(0+(in_buffer[2]<<1))-(0+(in_buffer[3]<<0)+(in_buffer[3]<<2)+(in_buffer[3]<<5)+(in_buffer[3]<<7))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2))+(0+(in_buffer[5]<<1)+(in_buffer[5]<<3)+(in_buffer[5]<<4)+(in_buffer[5]<<7))-(0+(in_buffer[6]<<0)+(in_buffer[6]<<2))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<4)+(in_buffer[7]<<5))+(0+(in_buffer[8]<<2)+(in_buffer[8]<<4)+(in_buffer[8]<<6))+(0-(in_buffer[9]<<1)-(in_buffer[9]<<3)+(in_buffer[9]<<5)+(in_buffer[9]<<6))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<4))+(0+(in_buffer[11]<<2)+(in_buffer[11]<<5)+(in_buffer[11]<<6))-(0-(in_buffer[12]<<2)+(in_buffer[12]<<6)+(in_buffer[12]<<7))+(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<1)+(in_buffer[14]<<2))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3))+(0-(in_buffer[16]<<0)+(in_buffer[16]<<3)+(in_buffer[16]<<4))+(0+(in_buffer[17]<<1)+(in_buffer[17]<<2)+(in_buffer[17]<<5))-(0+(in_buffer[18]<<0)-(in_buffer[18]<<3)+(in_buffer[18]<<7))+(0-(in_buffer[19]<<0)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<3)+(in_buffer[20]<<4))-(0+(in_buffer[21]<<0)+(in_buffer[21]<<1)+(in_buffer[21]<<4))-(0+(in_buffer[22]<<3)+(in_buffer[22]<<4))+(0+(in_buffer[23]<<3))-(0+(in_buffer[24]<<5))+(0+(in_buffer[25]<<3)+(in_buffer[25]<<6))+(0+(in_buffer[26]<<1)+(in_buffer[26]<<2)+(in_buffer[26]<<5))-(0+(in_buffer[27]<<0)+(in_buffer[27]<<2)+(in_buffer[27]<<5))-(0+(in_buffer[28]<<0)+(in_buffer[28]<<6))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<2)+(in_buffer[29]<<4)+(in_buffer[29]<<5))-(0-(in_buffer[30]<<0)-(in_buffer[30]<<3)+(in_buffer[30]<<6)+(in_buffer[30]<<7))+(0+(in_buffer[31]<<2))-(0+(in_buffer[32]<<2)+(in_buffer[32]<<5)+(in_buffer[32]<<7))+(0+(in_buffer[33]<<2)+(in_buffer[33]<<3))+(0+(in_buffer[34]<<3)+(in_buffer[34]<<5))+(0+(in_buffer[35]<<0)+(in_buffer[35]<<2)+(in_buffer[35]<<4)+(in_buffer[35]<<6))+(0-(in_buffer[36]<<1)+(in_buffer[36]<<4)+(in_buffer[36]<<6))+(0+(in_buffer[37]<<1)+(in_buffer[37]<<2)+(in_buffer[37]<<6))-(0-(in_buffer[38]<<0)-(in_buffer[38]<<3)+(in_buffer[38]<<5)+(in_buffer[38]<<6))+(0+(in_buffer[39]<<2)+(in_buffer[39]<<3)+(in_buffer[39]<<6))-(0+(in_buffer[40]<<1)+(in_buffer[40]<<3))+(0-(in_buffer[41]<<2)+(in_buffer[41]<<6))-(0+(in_buffer[42]<<0)+(in_buffer[42]<<2)+(in_buffer[42]<<3))-(0+(in_buffer[43]<<0)+(in_buffer[43]<<1)+(in_buffer[43]<<5)+(in_buffer[43]<<7))+(0+(in_buffer[44]<<0)+(in_buffer[44]<<2)+(in_buffer[44]<<4)+(in_buffer[44]<<5))+(0+(in_buffer[45]<<3)+(in_buffer[45]<<5))+(0+(in_buffer[46]<<0)+(in_buffer[46]<<3)+(in_buffer[46]<<5)+(in_buffer[46]<<6))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<2))+(0-(in_buffer[48]<<0)-(in_buffer[48]<<2)+(in_buffer[48]<<4)+(in_buffer[48]<<5))+(0+(in_buffer[49]<<0)+(in_buffer[49]<<1)+(in_buffer[49]<<4)+(in_buffer[49]<<5))+(0+(in_buffer[50]<<0)-(in_buffer[50]<<3)+(in_buffer[50]<<5)+(in_buffer[50]<<6))-(0+(in_buffer[51]<<3)+(in_buffer[51]<<5)+(in_buffer[51]<<7))-(0-(in_buffer[52]<<2)+(in_buffer[52]<<6)+(in_buffer[52]<<7))-(0+(in_buffer[53]<<0)-(in_buffer[53]<<3)+(in_buffer[53]<<7))-(0+(in_buffer[54]<<0)+(in_buffer[54]<<2)+(in_buffer[54]<<4))-(0-(in_buffer[55]<<1)+(in_buffer[55]<<7))-(0+(in_buffer[56]<<3)+(in_buffer[56]<<6))-(0+(in_buffer[57]<<0)+(in_buffer[57]<<1)+(in_buffer[57]<<4)+(in_buffer[57]<<5))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<3)+(in_buffer[58]<<4))-(0-(in_buffer[59]<<0)+(in_buffer[59]<<3))-(0+(in_buffer[60]<<2)+(in_buffer[60]<<4))+(0+(in_buffer[61]<<1)+(in_buffer[61]<<4)+(in_buffer[61]<<5))+(0+(in_buffer[62]<<0)+(in_buffer[62]<<1)+(in_buffer[62]<<6))-(0+(in_buffer[63]<<0)+(in_buffer[63]<<2)+(in_buffer[63]<<4)+(in_buffer[63]<<6)+(in_buffer[63]<<7));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight5;
assign in_buffer_weight5=0-(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<7))-(0+(in_buffer[2]<<3)+(in_buffer[2]<<5))+(0-(in_buffer[3]<<0)-(in_buffer[3]<<2)+(in_buffer[3]<<4)+(in_buffer[3]<<5))-(0+(in_buffer[4]<<0)+(in_buffer[4]<<2)-(in_buffer[4]<<5)+(in_buffer[4]<<8))-(0+(in_buffer[5]<<1)+(in_buffer[5]<<5))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<2)+(in_buffer[6]<<3))-(0+(in_buffer[7]<<0)-(in_buffer[7]<<2)+(in_buffer[7]<<5))+(0-(in_buffer[8]<<0)+(in_buffer[8]<<5)+(in_buffer[8]<<6))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<3)+(in_buffer[9]<<5)+(in_buffer[9]<<6))+(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)+(in_buffer[10]<<4))-(0-(in_buffer[11]<<0)-(in_buffer[11]<<3)+(in_buffer[11]<<6))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<3))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<2)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<2)+(in_buffer[14]<<3))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<1))+(0-(in_buffer[16]<<1)-(in_buffer[16]<<3)+(in_buffer[16]<<6))-(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4))-(0+(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<5))-(0-(in_buffer[19]<<3)+(in_buffer[19]<<5)+(in_buffer[19]<<6))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<3))+(0+(in_buffer[21]<<0)+(in_buffer[21]<<5))-(0+(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<4)+(in_buffer[22]<<5))+(0+(in_buffer[23]<<1)+(in_buffer[23]<<3)+(in_buffer[23]<<6))-(0-(in_buffer[24]<<1)+(in_buffer[24]<<4))+(0+(in_buffer[25]<<0)+(in_buffer[25]<<1)+(in_buffer[25]<<4))+(0-(in_buffer[26]<<0)+(in_buffer[26]<<3)+(in_buffer[26]<<5)+(in_buffer[26]<<6))+(0+(in_buffer[27]<<1)+(in_buffer[27]<<3)+(in_buffer[27]<<4))-(0-(in_buffer[28]<<0)+(in_buffer[28]<<2)+(in_buffer[28]<<3)+(in_buffer[28]<<7))-(0+(in_buffer[29]<<1)+(in_buffer[29]<<4)+(in_buffer[29]<<6))+(0-(in_buffer[30]<<1)+(in_buffer[30]<<7))+(0+(in_buffer[31]<<0))+(0+(in_buffer[32]<<4)+(in_buffer[32]<<5))+(0-(in_buffer[33]<<2)+(in_buffer[33]<<5))+(0+(in_buffer[35]<<2)+(in_buffer[35]<<5))-(0+(in_buffer[36]<<0)+(in_buffer[36]<<2))+(0-(in_buffer[37]<<0)-(in_buffer[37]<<3)+(in_buffer[37]<<6))+(0+(in_buffer[38]<<2))+(0-(in_buffer[39]<<1)+(in_buffer[39]<<3)+(in_buffer[39]<<4))-(0+(in_buffer[40]<<4))-(0+(in_buffer[41]<<0)+(in_buffer[41]<<3)+(in_buffer[41]<<4))-(0+(in_buffer[42]<<0)-(in_buffer[42]<<3)+(in_buffer[42]<<5)+(in_buffer[42]<<6))+(0+(in_buffer[43]<<2)+(in_buffer[43]<<5)+(in_buffer[43]<<6))-(0-(in_buffer[44]<<0)+(in_buffer[44]<<2)+(in_buffer[44]<<3))+(0-(in_buffer[45]<<0)+(in_buffer[45]<<2)+(in_buffer[45]<<3))-(0-(in_buffer[46]<<0)+(in_buffer[46]<<4)+(in_buffer[46]<<6))+(0+(in_buffer[47]<<1)+(in_buffer[47]<<3))+(0-(in_buffer[48]<<0)+(in_buffer[48]<<4))-(0-(in_buffer[49]<<0)+(in_buffer[49]<<3)+(in_buffer[49]<<5))+(0-(in_buffer[50]<<0)+(in_buffer[50]<<5))-(0-(in_buffer[51]<<0)+(in_buffer[51]<<4))+(0-(in_buffer[52]<<0)-(in_buffer[52]<<2)+(in_buffer[52]<<5)+(in_buffer[52]<<6))-(0+(in_buffer[53]<<1)+(in_buffer[53]<<4))-(0+(in_buffer[54]<<0)+(in_buffer[54]<<1)+(in_buffer[54]<<4)+(in_buffer[54]<<5))+(0+(in_buffer[55]<<2)+(in_buffer[55]<<3))+(0+(in_buffer[56]<<0)+(in_buffer[56]<<4)+(in_buffer[56]<<5))+(0-(in_buffer[57]<<2)+(in_buffer[57]<<5))-(0-(in_buffer[58]<<1)-(in_buffer[58]<<3)+(in_buffer[58]<<6))-(0+(in_buffer[59]<<3))-(0+(in_buffer[60]<<1)+(in_buffer[60]<<4))-(0+(in_buffer[61]<<6))+(0+(in_buffer[62]<<1)+(in_buffer[62]<<3))+(0-(in_buffer[63]<<0)+(in_buffer[63]<<2)+(in_buffer[63]<<3)+(in_buffer[63]<<6));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight6;
assign in_buffer_weight6=0+(0+(in_buffer[0]<<3))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<5))+(0+(in_buffer[2]<<4))+(0-(in_buffer[3]<<0)+(in_buffer[3]<<6))-(0-(in_buffer[4]<<0)+(in_buffer[4]<<2)+(in_buffer[4]<<3)+(in_buffer[4]<<7))+(0+(in_buffer[5]<<2)+(in_buffer[5]<<6))+(0-(in_buffer[6]<<0)+(in_buffer[6]<<4)+(in_buffer[6]<<5))-(0-(in_buffer[7]<<0)+(in_buffer[7]<<2)+(in_buffer[7]<<3))-(0-(in_buffer[8]<<1)-(in_buffer[8]<<3)+(in_buffer[8]<<6))+(0+(in_buffer[9]<<1)+(in_buffer[9]<<2))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<2)+(in_buffer[10]<<3))-(0+(in_buffer[11]<<3)+(in_buffer[11]<<5))+(0+(in_buffer[12]<<0)+(in_buffer[12]<<5))+(0-(in_buffer[13]<<0)-(in_buffer[13]<<2)+(in_buffer[13]<<4)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<2)+(in_buffer[14]<<3))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<4))-(0-(in_buffer[16]<<0)+(in_buffer[16]<<2)+(in_buffer[16]<<3)+(in_buffer[16]<<7))-(0+(in_buffer[17]<<0)-(in_buffer[17]<<2)+(in_buffer[17]<<6))+(0-(in_buffer[18]<<1)+(in_buffer[18]<<4)+(in_buffer[18]<<5))-(0-(in_buffer[19]<<1)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<0)+(in_buffer[20]<<2)+(in_buffer[20]<<3))+(0-(in_buffer[21]<<0)+(in_buffer[21]<<4))-(0-(in_buffer[22]<<0)-(in_buffer[22]<<2)+(in_buffer[22]<<6))-(0+(in_buffer[23]<<1)-(in_buffer[23]<<3)+(in_buffer[23]<<6))+(0+(in_buffer[24]<<0)+(in_buffer[24]<<3)+(in_buffer[24]<<5))-(0-(in_buffer[25]<<1)-(in_buffer[25]<<3)+(in_buffer[25]<<5)+(in_buffer[25]<<6))+(0+(in_buffer[26]<<3))+(0-(in_buffer[27]<<0)+(in_buffer[27]<<3)+(in_buffer[27]<<4))+(0+(in_buffer[28]<<0)+(in_buffer[28]<<2)+(in_buffer[28]<<5)+(in_buffer[28]<<6))-(0+(in_buffer[29]<<0)+(in_buffer[29]<<4)+(in_buffer[29]<<6))+(0-(in_buffer[30]<<1)+(in_buffer[30]<<4)+(in_buffer[30]<<7))-(0+(in_buffer[31]<<0)+(in_buffer[31]<<2))+(0-(in_buffer[32]<<0)+(in_buffer[32]<<7))+(0+(in_buffer[33]<<2)+(in_buffer[33]<<4)+(in_buffer[33]<<6))-(0+(in_buffer[35]<<0)+(in_buffer[35]<<1)-(in_buffer[35]<<4)+(in_buffer[35]<<7))-(0+(in_buffer[36]<<0)+(in_buffer[36]<<2)+(in_buffer[36]<<4)+(in_buffer[36]<<7)+(in_buffer[36]<<8))+(0+(in_buffer[37]<<0)+(in_buffer[37]<<4))-(0-(in_buffer[38]<<0)+(in_buffer[38]<<3))-(0+(in_buffer[39]<<2)+(in_buffer[39]<<7)+(in_buffer[39]<<8))-(0+(in_buffer[40]<<0)+(in_buffer[40]<<3))-(0+(in_buffer[41]<<2)+(in_buffer[41]<<5))-(0-(in_buffer[42]<<3)+(in_buffer[42]<<6))-(0+(in_buffer[43]<<1)+(in_buffer[43]<<4)+(in_buffer[43]<<6))+(0-(in_buffer[44]<<0)-(in_buffer[44]<<2)+(in_buffer[44]<<4)+(in_buffer[44]<<5))-(0-(in_buffer[45]<<2)+(in_buffer[45]<<4)+(in_buffer[45]<<5))+(0-(in_buffer[46]<<1)+(in_buffer[46]<<4)+(in_buffer[46]<<5))-(0-(in_buffer[47]<<0)+(in_buffer[47]<<3))-(0+(in_buffer[48]<<0)+(in_buffer[48]<<4)+(in_buffer[48]<<5))-(0-(in_buffer[49]<<0)+(in_buffer[49]<<3)+(in_buffer[49]<<7))-(0+(in_buffer[50]<<0)+(in_buffer[50]<<1))-(0+(in_buffer[51]<<0)+(in_buffer[51]<<2)+(in_buffer[51]<<6))-(0-(in_buffer[52]<<0)-(in_buffer[52]<<3)+(in_buffer[52]<<6))-(0+(in_buffer[53]<<3)+(in_buffer[53]<<6)+(in_buffer[53]<<7))+(0-(in_buffer[54]<<3)+(in_buffer[54]<<7))+(0-(in_buffer[55]<<1)+(in_buffer[55]<<4)+(in_buffer[55]<<6))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<4))+(0-(in_buffer[57]<<0)+(in_buffer[57]<<7))+(0+(in_buffer[58]<<1)+(in_buffer[58]<<4)+(in_buffer[58]<<5))-(0-(in_buffer[59]<<0)+(in_buffer[59]<<3))-(0+(in_buffer[60]<<0)+(in_buffer[60]<<2)+(in_buffer[60]<<6))-(0+(in_buffer[61]<<6))+(0+(in_buffer[62]<<1)+(in_buffer[62]<<3)+(in_buffer[62]<<5))+(0-(in_buffer[63]<<0)+(in_buffer[63]<<2)+(in_buffer[63]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight7;
assign in_buffer_weight7=0-(0-(in_buffer[0]<<0)+(in_buffer[0]<<3))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<1)+(in_buffer[1]<<4)+(in_buffer[1]<<5))+(0-(in_buffer[2]<<1)+(in_buffer[2]<<4))-(0+(in_buffer[3]<<1)-(in_buffer[3]<<4)+(in_buffer[3]<<7))+(0+(in_buffer[4]<<0)-(in_buffer[4]<<3)+(in_buffer[4]<<6))-(0+(in_buffer[5]<<0)+(in_buffer[5]<<3)+(in_buffer[5]<<6))-(0-(in_buffer[6]<<1)+(in_buffer[6]<<4)+(in_buffer[6]<<6))-(0-(in_buffer[7]<<4)+(in_buffer[7]<<7))-(0-(in_buffer[8]<<0)+(in_buffer[8]<<5)+(in_buffer[8]<<7))-(0+(in_buffer[9]<<2))-(0+(in_buffer[10]<<0)+(in_buffer[10]<<1)+(in_buffer[10]<<4))+(0-(in_buffer[11]<<0)+(in_buffer[11]<<4))+(0-(in_buffer[12]<<2)+(in_buffer[12]<<7))-(0+(in_buffer[13]<<4)+(in_buffer[13]<<5))-(0+(in_buffer[14]<<3))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<2)+(in_buffer[15]<<3))+(0+(in_buffer[16]<<4)+(in_buffer[16]<<5))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4))-(0-(in_buffer[18]<<0)+(in_buffer[18]<<5))+(0+(in_buffer[19]<<0)+(in_buffer[19]<<3)+(in_buffer[19]<<5))+(0+(in_buffer[20]<<2))+(0+(in_buffer[22]<<1)+(in_buffer[22]<<3)+(in_buffer[22]<<5))+(0+(in_buffer[23]<<2)+(in_buffer[23]<<4))-(0+(in_buffer[24]<<1)+(in_buffer[24]<<3))-(0+(in_buffer[25]<<1)+(in_buffer[25]<<2))+(0+(in_buffer[26]<<2)+(in_buffer[26]<<6))+(0+(in_buffer[27]<<1)+(in_buffer[27]<<3))-(0-(in_buffer[28]<<0)+(in_buffer[28]<<3))+(0+(in_buffer[29]<<0)+(in_buffer[29]<<3)+(in_buffer[29]<<5)+(in_buffer[29]<<6))-(0+(in_buffer[30]<<2)+(in_buffer[30]<<7))-(0+(in_buffer[31]<<1)+(in_buffer[31]<<3))-(0-(in_buffer[32]<<0)-(in_buffer[32]<<2)+(in_buffer[32]<<5)+(in_buffer[32]<<6))-(0-(in_buffer[33]<<0)-(in_buffer[33]<<2)+(in_buffer[33]<<4)+(in_buffer[33]<<5))-(0-(in_buffer[34]<<2)+(in_buffer[34]<<5)+(in_buffer[34]<<6))+(0-(in_buffer[35]<<1)+(in_buffer[35]<<4)+(in_buffer[35]<<6))+(0+(in_buffer[36]<<0)+(in_buffer[36]<<1)+(in_buffer[36]<<4)+(in_buffer[36]<<5))-(0+(in_buffer[37]<<1)-(in_buffer[37]<<3)+(in_buffer[37]<<6))+(0+(in_buffer[38]<<3)+(in_buffer[38]<<4))-(0+(in_buffer[39]<<0)+(in_buffer[39]<<4))-(0+(in_buffer[40]<<0)+(in_buffer[40]<<3))+(0+(in_buffer[41]<<0)-(in_buffer[41]<<3)+(in_buffer[41]<<6))+(0-(in_buffer[42]<<1)+(in_buffer[42]<<7))-(0+(in_buffer[43]<<2)+(in_buffer[43]<<3)+(in_buffer[43]<<6))-(0+(in_buffer[44]<<0)+(in_buffer[44]<<2)+(in_buffer[44]<<5))-(0-(in_buffer[45]<<1)+(in_buffer[45]<<7))-(0+(in_buffer[46]<<2)+(in_buffer[46]<<4))+(0+(in_buffer[47]<<0)+(in_buffer[47]<<2))+(0+(in_buffer[48]<<2)+(in_buffer[48]<<6))+(0+(in_buffer[49]<<0)+(in_buffer[49]<<4)+(in_buffer[49]<<5))+(0+(in_buffer[50]<<2)+(in_buffer[50]<<4))+(0-(in_buffer[51]<<0)+(in_buffer[51]<<4))-(0+(in_buffer[52]<<1)+(in_buffer[52]<<5))+(0+(in_buffer[53]<<0)+(in_buffer[53]<<2)+(in_buffer[53]<<3)+(in_buffer[53]<<6))+(0-(in_buffer[54]<<0)+(in_buffer[54]<<3)+(in_buffer[54]<<4))-(0-(in_buffer[55]<<0)+(in_buffer[55]<<4))-(0+(in_buffer[56]<<0)+(in_buffer[56]<<2)+(in_buffer[56]<<4))+(0+(in_buffer[57]<<0)+(in_buffer[57]<<4))+(0+(in_buffer[58]<<1)+(in_buffer[58]<<2)+(in_buffer[58]<<6))+(0-(in_buffer[60]<<0)-(in_buffer[60]<<2)+(in_buffer[60]<<5))+(0-(in_buffer[61]<<1)+(in_buffer[61]<<5))+(0+(in_buffer[62]<<0)+(in_buffer[62]<<1))-(0+(in_buffer[63]<<2)+(in_buffer[63]<<5));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight8;
assign in_buffer_weight8=0+(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3))-(0+(in_buffer[1]<<0)+(in_buffer[1]<<1)+(in_buffer[1]<<4))+(0+(in_buffer[2]<<0)+(in_buffer[2]<<4))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<2))-(0-(in_buffer[4]<<3)+(in_buffer[4]<<6))-(0-(in_buffer[5]<<1)+(in_buffer[5]<<3)+(in_buffer[5]<<4))+(0+(in_buffer[6]<<0)-(in_buffer[6]<<3)+(in_buffer[6]<<6))+(0+(in_buffer[7]<<1)+(in_buffer[7]<<2)+(in_buffer[7]<<5))+(0-(in_buffer[8]<<1)+(in_buffer[8]<<4)+(in_buffer[8]<<5))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<6))+(0+(in_buffer[10]<<4))-(0+(in_buffer[11]<<0)-(in_buffer[11]<<4)+(in_buffer[11]<<7))-(0+(in_buffer[12]<<0)-(in_buffer[12]<<2)+(in_buffer[12]<<4)+(in_buffer[12]<<5))+(0-(in_buffer[13]<<0)+(in_buffer[13]<<5))-(0-(in_buffer[14]<<0)+(in_buffer[14]<<3))+(0-(in_buffer[15]<<0)+(in_buffer[15]<<3))-(0+(in_buffer[16]<<1)+(in_buffer[16]<<2)+(in_buffer[16]<<5))-(0+(in_buffer[17]<<1)+(in_buffer[17]<<2))-(0+(in_buffer[18]<<0)-(in_buffer[18]<<2)+(in_buffer[18]<<5))-(0+(in_buffer[19]<<0)+(in_buffer[19]<<3)+(in_buffer[19]<<5)+(in_buffer[19]<<8))+(0+(in_buffer[20]<<1)+(in_buffer[20]<<2))+(0+(in_buffer[21]<<5))+(0+(in_buffer[22]<<3)+(in_buffer[22]<<5))-(0-(in_buffer[23]<<0)+(in_buffer[23]<<6))+(0+(in_buffer[24]<<2))-(0-(in_buffer[25]<<0)+(in_buffer[25]<<4))-(0-(in_buffer[26]<<0)+(in_buffer[26]<<3)+(in_buffer[26]<<5))+(0-(in_buffer[27]<<2)+(in_buffer[27]<<5))+(0+(in_buffer[28]<<4))+(0+(in_buffer[29]<<1))-(0+(in_buffer[30]<<2)+(in_buffer[30]<<5))-(0-(in_buffer[31]<<0)+(in_buffer[31]<<3))+(0+(in_buffer[32]<<4)+(in_buffer[32]<<5))-(0+(in_buffer[33]<<0)+(in_buffer[33]<<1)+(in_buffer[33]<<4))-(0+(in_buffer[34]<<1)+(in_buffer[34]<<2)+(in_buffer[34]<<5)+(in_buffer[34]<<6))-(0+(in_buffer[35]<<0)+(in_buffer[35]<<2)+(in_buffer[35]<<3))+(0+(in_buffer[36]<<1)+(in_buffer[36]<<3)+(in_buffer[36]<<5))+(0-(in_buffer[37]<<0)+(in_buffer[37]<<6))+(0+(in_buffer[38]<<2)+(in_buffer[38]<<5)+(in_buffer[38]<<6))-(0+(in_buffer[39]<<1)+(in_buffer[39]<<2)+(in_buffer[39]<<7))+(0+(in_buffer[40]<<1)+(in_buffer[40]<<2))-(0+(in_buffer[41]<<1)+(in_buffer[41]<<6))-(0+(in_buffer[42]<<0)-(in_buffer[42]<<3)+(in_buffer[42]<<6))-(0+(in_buffer[43]<<0)+(in_buffer[43]<<3)+(in_buffer[43]<<4))-(0+(in_buffer[44]<<3)+(in_buffer[44]<<4))+(0-(in_buffer[45]<<2)+(in_buffer[45]<<5))-(0-(in_buffer[46]<<1)+(in_buffer[46]<<5)+(in_buffer[46]<<6))-(0+(in_buffer[48]<<0)+(in_buffer[48]<<2))+(0+(in_buffer[49]<<2)+(in_buffer[49]<<4))-(0+(in_buffer[50]<<1)+(in_buffer[50]<<3))+(0-(in_buffer[51]<<1)+(in_buffer[51]<<3)+(in_buffer[51]<<4))+(0-(in_buffer[52]<<1)+(in_buffer[52]<<3)+(in_buffer[52]<<4))-(0+(in_buffer[53]<<0)-(in_buffer[53]<<3)+(in_buffer[53]<<6))+(0+(in_buffer[54]<<1)+(in_buffer[54]<<3))-(0+(in_buffer[55]<<0)+(in_buffer[55]<<1)+(in_buffer[55]<<4)+(in_buffer[55]<<5))-(0+(in_buffer[56]<<1)+(in_buffer[56]<<3))-(0+(in_buffer[57]<<0)+(in_buffer[57]<<3)+(in_buffer[57]<<4))-(0+(in_buffer[58]<<1)+(in_buffer[58]<<5)+(in_buffer[58]<<6))+(0+(in_buffer[59]<<1))+(0-(in_buffer[60]<<0)-(in_buffer[60]<<2)+(in_buffer[60]<<5))+(0+(in_buffer[61]<<0)+(in_buffer[61]<<2)+(in_buffer[61]<<3))+(0+(in_buffer[62]<<0)+(in_buffer[62]<<3)+(in_buffer[62]<<4))+(0+(in_buffer[63]<<0)+(in_buffer[63]<<3));
wire signed  [DATA_WIDTH-1:0]   in_buffer_weight9;
assign in_buffer_weight9=0-(0+(in_buffer[0]<<0)+(in_buffer[0]<<2)+(in_buffer[0]<<3))+(0+(in_buffer[1]<<0)+(in_buffer[1]<<2)+(in_buffer[1]<<3))+(0+(in_buffer[3]<<1)+(in_buffer[3]<<2)+(in_buffer[3]<<5))+(0-(in_buffer[4]<<0)+(in_buffer[4]<<6))-(0+(in_buffer[5]<<0)-(in_buffer[5]<<2)+(in_buffer[5]<<6)+(in_buffer[5]<<7))+(0+(in_buffer[6]<<0)+(in_buffer[6]<<1))+(0-(in_buffer[7]<<0)-(in_buffer[7]<<2)+(in_buffer[7]<<5))+(0+(in_buffer[8]<<4)+(in_buffer[8]<<5))-(0+(in_buffer[9]<<0)+(in_buffer[9]<<1)+(in_buffer[9]<<6))-(0+(in_buffer[10]<<0)-(in_buffer[10]<<2)+(in_buffer[10]<<5))-(0-(in_buffer[11]<<1)+(in_buffer[11]<<3)+(in_buffer[11]<<4))-(0-(in_buffer[12]<<1)+(in_buffer[12]<<4)+(in_buffer[12]<<6))-(0+(in_buffer[13]<<0)+(in_buffer[13]<<5))+(0+(in_buffer[14]<<2))-(0+(in_buffer[15]<<0)+(in_buffer[15]<<1))+(0+(in_buffer[16]<<1)+(in_buffer[16]<<3)+(in_buffer[16]<<4))+(0+(in_buffer[17]<<0)+(in_buffer[17]<<1)+(in_buffer[17]<<4)+(in_buffer[17]<<5))+(0+(in_buffer[18]<<3)+(in_buffer[18]<<4))+(0+(in_buffer[19]<<2)+(in_buffer[19]<<5))+(0-(in_buffer[20]<<2)+(in_buffer[20]<<5))+(0+(in_buffer[21]<<4)+(in_buffer[21]<<5))-(0+(in_buffer[22]<<0)+(in_buffer[22]<<3)+(in_buffer[22]<<6))+(0+(in_buffer[23]<<4)+(in_buffer[23]<<6))-(0+(in_buffer[24]<<1)+(in_buffer[24]<<3)+(in_buffer[24]<<5))-(0-(in_buffer[25]<<0)+(in_buffer[25]<<8))-(0-(in_buffer[26]<<2)+(in_buffer[26]<<6))-(0+(in_buffer[28]<<4)+(in_buffer[28]<<6))+(0+(in_buffer[29]<<2)+(in_buffer[29]<<4))-(0+(in_buffer[30]<<0)+(in_buffer[30]<<4)+(in_buffer[30]<<5))+(0+(in_buffer[31]<<0))-(0+(in_buffer[32]<<0)+(in_buffer[32]<<1)+(in_buffer[32]<<5))+(0+(in_buffer[33]<<1)+(in_buffer[33]<<2)+(in_buffer[33]<<6))+(0-(in_buffer[34]<<0)-(in_buffer[34]<<3)+(in_buffer[34]<<7))+(0+(in_buffer[35]<<4)+(in_buffer[35]<<5))+(0+(in_buffer[36]<<1)+(in_buffer[36]<<3))+(0+(in_buffer[37]<<4))-(0+(in_buffer[38]<<0)+(in_buffer[38]<<4)+(in_buffer[38]<<6))+(0-(in_buffer[39]<<0)+(in_buffer[39]<<6))-(0+(in_buffer[40]<<1)+(in_buffer[40]<<2))+(0+(in_buffer[41]<<0)+(in_buffer[41]<<4))+(0+(in_buffer[42]<<0)+(in_buffer[42]<<2))+(0+(in_buffer[43]<<0))+(0+(in_buffer[44]<<4))-(0+(in_buffer[45]<<0)+(in_buffer[45]<<3))-(0-(in_buffer[46]<<1)-(in_buffer[46]<<4)+(in_buffer[46]<<6)+(in_buffer[46]<<7))-(0+(in_buffer[47]<<2)+(in_buffer[47]<<3))+(0+(in_buffer[48]<<0)-(in_buffer[48]<<2)+(in_buffer[48]<<5))+(0-(in_buffer[49]<<2)+(in_buffer[49]<<5))-(0+(in_buffer[50]<<0)+(in_buffer[50]<<6))-(0+(in_buffer[51]<<1)+(in_buffer[51]<<4))-(0-(in_buffer[52]<<0)+(in_buffer[52]<<4)+(in_buffer[52]<<6))-(0-(in_buffer[53]<<0)+(in_buffer[53]<<3)+(in_buffer[53]<<5)+(in_buffer[53]<<6))-(0+(in_buffer[54]<<2)+(in_buffer[54]<<3)+(in_buffer[54]<<6))+(0+(in_buffer[55]<<0)+(in_buffer[55]<<1))-(0+(in_buffer[57]<<1)-(in_buffer[57]<<3)-(in_buffer[57]<<5)+(in_buffer[57]<<8))-(0+(in_buffer[58]<<0)+(in_buffer[58]<<2)+(in_buffer[58]<<5)+(in_buffer[58]<<6))-(0+(in_buffer[59]<<2))+(0-(in_buffer[60]<<0)-(in_buffer[60]<<2)+(in_buffer[60]<<4)+(in_buffer[60]<<5))+(0+(in_buffer[61]<<1)+(in_buffer[61]<<3)+(in_buffer[61]<<5))-(0-(in_buffer[62]<<0)+(in_buffer[62]<<5)+(in_buffer[62]<<7))+(0+(in_buffer[63]<<0)+(in_buffer[63]<<4));
wire signed [DATA_WIDTH-1:0]   weight_bias0;
wire signed [DATA_WIDTH-1:0]   weight_bias1;
wire signed [DATA_WIDTH-1:0]   weight_bias2;
wire signed [DATA_WIDTH-1:0]   weight_bias3;
wire signed [DATA_WIDTH-1:0]   weight_bias4;
wire signed [DATA_WIDTH-1:0]   weight_bias5;
wire signed [DATA_WIDTH-1:0]   weight_bias6;
wire signed [DATA_WIDTH-1:0]   weight_bias7;
wire signed [DATA_WIDTH-1:0]   weight_bias8;
wire signed [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias0=in_buffer_weight0+(-49);
assign weight_bias1=in_buffer_weight1+(-1);
assign weight_bias2=in_buffer_weight2+(51);
assign weight_bias3=in_buffer_weight3+(-30);
assign weight_bias4=in_buffer_weight4+(-29);
assign weight_bias5=in_buffer_weight5+(27);
assign weight_bias6=in_buffer_weight6+(11);
assign weight_bias7=in_buffer_weight7+(-21);
assign weight_bias8=in_buffer_weight8+(3);
assign weight_bias9=in_buffer_weight9+(29);
assign layer_out={weight_bias9,weight_bias8,weight_bias7,weight_bias6,weight_bias5,weight_bias4,weight_bias3,weight_bias2,weight_bias1,weight_bias0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule