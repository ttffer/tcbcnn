//version 1 constant in Verilog
module con1
    #(
        parameter   OUTPUT_BIT  =   19,
                    OUTPUT_NODE =   100,
                    DATA_WIDTH  =   19,
                    IMG_SZ    =   11*11
)
(
    input   clk,
    input   rst,
    input   [IMG_SZ*8-1:0]   img,
    input   valid,
    output  reg ready,
    output [OUTPUT_BIT*OUTPUT_NODE-1:0] layer_out
);

reg    signed [8-1:0]  in_buffer[0:IMG_SZ-1];
genvar j;
generate
for(j=0;j<IMG_SZ;j=j+1) 
    begin:init_block
        always@(posedge clk)
            begin
                if(rst)
                    begin
                        in_buffer[j]<=0;
                    end
                else
                    begin
                        in_buffer[j]<=img[j*8+7:j*8+0];
                    end
            end
    end
endgenerate
//wire declatation
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight0;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight1;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight2;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight3;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight4;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight5;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight6;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight7;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight8;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight9;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight10;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight11;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight12;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight13;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight14;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight15;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight16;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight17;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight18;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight19;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight20;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight21;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight22;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight23;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight24;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight25;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight26;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight27;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight28;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight29;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight30;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight31;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight32;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight33;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight34;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight35;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight36;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight37;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight38;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight39;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight40;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight41;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight42;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight43;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight44;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight45;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight46;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight47;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight48;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight49;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight50;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight51;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight52;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight53;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight54;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight55;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight56;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight57;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight58;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight59;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight60;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight61;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight62;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight63;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight64;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight65;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight66;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight67;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight68;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight69;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight70;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight71;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight72;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight73;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight74;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight75;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight76;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight77;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight78;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight79;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight80;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight81;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight82;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight83;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight84;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight85;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight86;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight87;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight88;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight89;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight90;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight91;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight92;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight93;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight94;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight95;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight96;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight97;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight98;
wire signed    [DATA_WIDTH-1:0]   in_buffer_weight99;
assign in_buffer_weight0=297*in_buffer[0]+262*in_buffer[1]+255*in_buffer[11]+308*in_buffer[12];
assign in_buffer_weight1=297*in_buffer[1]+262*in_buffer[2]+255*in_buffer[12]+308*in_buffer[13];
assign in_buffer_weight2=297*in_buffer[2]+262*in_buffer[3]+255*in_buffer[13]+308*in_buffer[14];
assign in_buffer_weight3=297*in_buffer[3]+262*in_buffer[4]+255*in_buffer[14]+308*in_buffer[15];
assign in_buffer_weight4=297*in_buffer[4]+262*in_buffer[5]+255*in_buffer[15]+308*in_buffer[16];
assign in_buffer_weight5=297*in_buffer[5]+262*in_buffer[6]+255*in_buffer[16]+308*in_buffer[17];
assign in_buffer_weight6=297*in_buffer[6]+262*in_buffer[7]+255*in_buffer[17]+308*in_buffer[18];
assign in_buffer_weight7=297*in_buffer[7]+262*in_buffer[8]+255*in_buffer[18]+308*in_buffer[19];
assign in_buffer_weight8=297*in_buffer[8]+262*in_buffer[9]+255*in_buffer[19]+308*in_buffer[20];
assign in_buffer_weight9=297*in_buffer[9]+262*in_buffer[10]+255*in_buffer[20]+308*in_buffer[21];
assign in_buffer_weight10=297*in_buffer[11]+262*in_buffer[12]+255*in_buffer[22]+308*in_buffer[23];
assign in_buffer_weight11=297*in_buffer[12]+262*in_buffer[13]+255*in_buffer[23]+308*in_buffer[24];
assign in_buffer_weight12=297*in_buffer[13]+262*in_buffer[14]+255*in_buffer[24]+308*in_buffer[25];
assign in_buffer_weight13=297*in_buffer[14]+262*in_buffer[15]+255*in_buffer[25]+308*in_buffer[26];
assign in_buffer_weight14=297*in_buffer[15]+262*in_buffer[16]+255*in_buffer[26]+308*in_buffer[27];
assign in_buffer_weight15=297*in_buffer[16]+262*in_buffer[17]+255*in_buffer[27]+308*in_buffer[28];
assign in_buffer_weight16=297*in_buffer[17]+262*in_buffer[18]+255*in_buffer[28]+308*in_buffer[29];
assign in_buffer_weight17=297*in_buffer[18]+262*in_buffer[19]+255*in_buffer[29]+308*in_buffer[30];
assign in_buffer_weight18=297*in_buffer[19]+262*in_buffer[20]+255*in_buffer[30]+308*in_buffer[31];
assign in_buffer_weight19=297*in_buffer[20]+262*in_buffer[21]+255*in_buffer[31]+308*in_buffer[32];
assign in_buffer_weight20=297*in_buffer[22]+262*in_buffer[23]+255*in_buffer[33]+308*in_buffer[34];
assign in_buffer_weight21=297*in_buffer[23]+262*in_buffer[24]+255*in_buffer[34]+308*in_buffer[35];
assign in_buffer_weight22=297*in_buffer[24]+262*in_buffer[25]+255*in_buffer[35]+308*in_buffer[36];
assign in_buffer_weight23=297*in_buffer[25]+262*in_buffer[26]+255*in_buffer[36]+308*in_buffer[37];
assign in_buffer_weight24=297*in_buffer[26]+262*in_buffer[27]+255*in_buffer[37]+308*in_buffer[38];
assign in_buffer_weight25=297*in_buffer[27]+262*in_buffer[28]+255*in_buffer[38]+308*in_buffer[39];
assign in_buffer_weight26=297*in_buffer[28]+262*in_buffer[29]+255*in_buffer[39]+308*in_buffer[40];
assign in_buffer_weight27=297*in_buffer[29]+262*in_buffer[30]+255*in_buffer[40]+308*in_buffer[41];
assign in_buffer_weight28=297*in_buffer[30]+262*in_buffer[31]+255*in_buffer[41]+308*in_buffer[42];
assign in_buffer_weight29=297*in_buffer[31]+262*in_buffer[32]+255*in_buffer[42]+308*in_buffer[43];
assign in_buffer_weight30=297*in_buffer[33]+262*in_buffer[34]+255*in_buffer[44]+308*in_buffer[45];
assign in_buffer_weight31=297*in_buffer[34]+262*in_buffer[35]+255*in_buffer[45]+308*in_buffer[46];
assign in_buffer_weight32=297*in_buffer[35]+262*in_buffer[36]+255*in_buffer[46]+308*in_buffer[47];
assign in_buffer_weight33=297*in_buffer[36]+262*in_buffer[37]+255*in_buffer[47]+308*in_buffer[48];
assign in_buffer_weight34=297*in_buffer[37]+262*in_buffer[38]+255*in_buffer[48]+308*in_buffer[49];
assign in_buffer_weight35=297*in_buffer[38]+262*in_buffer[39]+255*in_buffer[49]+308*in_buffer[50];
assign in_buffer_weight36=297*in_buffer[39]+262*in_buffer[40]+255*in_buffer[50]+308*in_buffer[51];
assign in_buffer_weight37=297*in_buffer[40]+262*in_buffer[41]+255*in_buffer[51]+308*in_buffer[52];
assign in_buffer_weight38=297*in_buffer[41]+262*in_buffer[42]+255*in_buffer[52]+308*in_buffer[53];
assign in_buffer_weight39=297*in_buffer[42]+262*in_buffer[43]+255*in_buffer[53]+308*in_buffer[54];
assign in_buffer_weight40=297*in_buffer[44]+262*in_buffer[45]+255*in_buffer[55]+308*in_buffer[56];
assign in_buffer_weight41=297*in_buffer[45]+262*in_buffer[46]+255*in_buffer[56]+308*in_buffer[57];
assign in_buffer_weight42=297*in_buffer[46]+262*in_buffer[47]+255*in_buffer[57]+308*in_buffer[58];
assign in_buffer_weight43=297*in_buffer[47]+262*in_buffer[48]+255*in_buffer[58]+308*in_buffer[59];
assign in_buffer_weight44=297*in_buffer[48]+262*in_buffer[49]+255*in_buffer[59]+308*in_buffer[60];
assign in_buffer_weight45=297*in_buffer[49]+262*in_buffer[50]+255*in_buffer[60]+308*in_buffer[61];
assign in_buffer_weight46=297*in_buffer[50]+262*in_buffer[51]+255*in_buffer[61]+308*in_buffer[62];
assign in_buffer_weight47=297*in_buffer[51]+262*in_buffer[52]+255*in_buffer[62]+308*in_buffer[63];
assign in_buffer_weight48=297*in_buffer[52]+262*in_buffer[53]+255*in_buffer[63]+308*in_buffer[64];
assign in_buffer_weight49=297*in_buffer[53]+262*in_buffer[54]+255*in_buffer[64]+308*in_buffer[65];
assign in_buffer_weight50=297*in_buffer[55]+262*in_buffer[56]+255*in_buffer[66]+308*in_buffer[67];
assign in_buffer_weight51=297*in_buffer[56]+262*in_buffer[57]+255*in_buffer[67]+308*in_buffer[68];
assign in_buffer_weight52=297*in_buffer[57]+262*in_buffer[58]+255*in_buffer[68]+308*in_buffer[69];
assign in_buffer_weight53=297*in_buffer[58]+262*in_buffer[59]+255*in_buffer[69]+308*in_buffer[70];
assign in_buffer_weight54=297*in_buffer[59]+262*in_buffer[60]+255*in_buffer[70]+308*in_buffer[71];
assign in_buffer_weight55=297*in_buffer[60]+262*in_buffer[61]+255*in_buffer[71]+308*in_buffer[72];
assign in_buffer_weight56=297*in_buffer[61]+262*in_buffer[62]+255*in_buffer[72]+308*in_buffer[73];
assign in_buffer_weight57=297*in_buffer[62]+262*in_buffer[63]+255*in_buffer[73]+308*in_buffer[74];
assign in_buffer_weight58=297*in_buffer[63]+262*in_buffer[64]+255*in_buffer[74]+308*in_buffer[75];
assign in_buffer_weight59=297*in_buffer[64]+262*in_buffer[65]+255*in_buffer[75]+308*in_buffer[76];
assign in_buffer_weight60=297*in_buffer[66]+262*in_buffer[67]+255*in_buffer[77]+308*in_buffer[78];
assign in_buffer_weight61=297*in_buffer[67]+262*in_buffer[68]+255*in_buffer[78]+308*in_buffer[79];
assign in_buffer_weight62=297*in_buffer[68]+262*in_buffer[69]+255*in_buffer[79]+308*in_buffer[80];
assign in_buffer_weight63=297*in_buffer[69]+262*in_buffer[70]+255*in_buffer[80]+308*in_buffer[81];
assign in_buffer_weight64=297*in_buffer[70]+262*in_buffer[71]+255*in_buffer[81]+308*in_buffer[82];
assign in_buffer_weight65=297*in_buffer[71]+262*in_buffer[72]+255*in_buffer[82]+308*in_buffer[83];
assign in_buffer_weight66=297*in_buffer[72]+262*in_buffer[73]+255*in_buffer[83]+308*in_buffer[84];
assign in_buffer_weight67=297*in_buffer[73]+262*in_buffer[74]+255*in_buffer[84]+308*in_buffer[85];
assign in_buffer_weight68=297*in_buffer[74]+262*in_buffer[75]+255*in_buffer[85]+308*in_buffer[86];
assign in_buffer_weight69=297*in_buffer[75]+262*in_buffer[76]+255*in_buffer[86]+308*in_buffer[87];
assign in_buffer_weight70=297*in_buffer[77]+262*in_buffer[78]+255*in_buffer[88]+308*in_buffer[89];
assign in_buffer_weight71=297*in_buffer[78]+262*in_buffer[79]+255*in_buffer[89]+308*in_buffer[90];
assign in_buffer_weight72=297*in_buffer[79]+262*in_buffer[80]+255*in_buffer[90]+308*in_buffer[91];
assign in_buffer_weight73=297*in_buffer[80]+262*in_buffer[81]+255*in_buffer[91]+308*in_buffer[92];
assign in_buffer_weight74=297*in_buffer[81]+262*in_buffer[82]+255*in_buffer[92]+308*in_buffer[93];
assign in_buffer_weight75=297*in_buffer[82]+262*in_buffer[83]+255*in_buffer[93]+308*in_buffer[94];
assign in_buffer_weight76=297*in_buffer[83]+262*in_buffer[84]+255*in_buffer[94]+308*in_buffer[95];
assign in_buffer_weight77=297*in_buffer[84]+262*in_buffer[85]+255*in_buffer[95]+308*in_buffer[96];
assign in_buffer_weight78=297*in_buffer[85]+262*in_buffer[86]+255*in_buffer[96]+308*in_buffer[97];
assign in_buffer_weight79=297*in_buffer[86]+262*in_buffer[87]+255*in_buffer[97]+308*in_buffer[98];
assign in_buffer_weight80=297*in_buffer[88]+262*in_buffer[89]+255*in_buffer[99]+308*in_buffer[100];
assign in_buffer_weight81=297*in_buffer[89]+262*in_buffer[90]+255*in_buffer[100]+308*in_buffer[101];
assign in_buffer_weight82=297*in_buffer[90]+262*in_buffer[91]+255*in_buffer[101]+308*in_buffer[102];
assign in_buffer_weight83=297*in_buffer[91]+262*in_buffer[92]+255*in_buffer[102]+308*in_buffer[103];
assign in_buffer_weight84=297*in_buffer[92]+262*in_buffer[93]+255*in_buffer[103]+308*in_buffer[104];
assign in_buffer_weight85=297*in_buffer[93]+262*in_buffer[94]+255*in_buffer[104]+308*in_buffer[105];
assign in_buffer_weight86=297*in_buffer[94]+262*in_buffer[95]+255*in_buffer[105]+308*in_buffer[106];
assign in_buffer_weight87=297*in_buffer[95]+262*in_buffer[96]+255*in_buffer[106]+308*in_buffer[107];
assign in_buffer_weight88=297*in_buffer[96]+262*in_buffer[97]+255*in_buffer[107]+308*in_buffer[108];
assign in_buffer_weight89=297*in_buffer[97]+262*in_buffer[98]+255*in_buffer[108]+308*in_buffer[109];
assign in_buffer_weight90=297*in_buffer[99]+262*in_buffer[100]+255*in_buffer[110]+308*in_buffer[111];
assign in_buffer_weight91=297*in_buffer[100]+262*in_buffer[101]+255*in_buffer[111]+308*in_buffer[112];
assign in_buffer_weight92=297*in_buffer[101]+262*in_buffer[102]+255*in_buffer[112]+308*in_buffer[113];
assign in_buffer_weight93=297*in_buffer[102]+262*in_buffer[103]+255*in_buffer[113]+308*in_buffer[114];
assign in_buffer_weight94=297*in_buffer[103]+262*in_buffer[104]+255*in_buffer[114]+308*in_buffer[115];
assign in_buffer_weight95=297*in_buffer[104]+262*in_buffer[105]+255*in_buffer[115]+308*in_buffer[116];
assign in_buffer_weight96=297*in_buffer[105]+262*in_buffer[106]+255*in_buffer[116]+308*in_buffer[117];
assign in_buffer_weight97=297*in_buffer[106]+262*in_buffer[107]+255*in_buffer[117]+308*in_buffer[118];
assign in_buffer_weight98=297*in_buffer[107]+262*in_buffer[108]+255*in_buffer[118]+308*in_buffer[119];
assign in_buffer_weight99=297*in_buffer[108]+262*in_buffer[109]+255*in_buffer[119]+308*in_buffer[120];
wire signed    [DATA_WIDTH-1:0]   weight_bias0;
assign weight_bias0= in_buffer_weight0+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias1;
assign weight_bias1= in_buffer_weight1+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias2;
assign weight_bias2= in_buffer_weight2+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias3;
assign weight_bias3= in_buffer_weight3+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias4;
assign weight_bias4= in_buffer_weight4+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias5;
assign weight_bias5= in_buffer_weight5+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias6;
assign weight_bias6= in_buffer_weight6+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias7;
assign weight_bias7= in_buffer_weight7+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias8;
assign weight_bias8= in_buffer_weight8+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias9;
assign weight_bias9= in_buffer_weight9+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias10;
assign weight_bias10= in_buffer_weight10+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias11;
assign weight_bias11= in_buffer_weight11+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias12;
assign weight_bias12= in_buffer_weight12+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias13;
assign weight_bias13= in_buffer_weight13+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias14;
assign weight_bias14= in_buffer_weight14+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias15;
assign weight_bias15= in_buffer_weight15+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias16;
assign weight_bias16= in_buffer_weight16+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias17;
assign weight_bias17= in_buffer_weight17+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias18;
assign weight_bias18= in_buffer_weight18+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias19;
assign weight_bias19= in_buffer_weight19+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias20;
assign weight_bias20= in_buffer_weight20+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias21;
assign weight_bias21= in_buffer_weight21+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias22;
assign weight_bias22= in_buffer_weight22+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias23;
assign weight_bias23= in_buffer_weight23+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias24;
assign weight_bias24= in_buffer_weight24+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias25;
assign weight_bias25= in_buffer_weight25+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias26;
assign weight_bias26= in_buffer_weight26+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias27;
assign weight_bias27= in_buffer_weight27+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias28;
assign weight_bias28= in_buffer_weight28+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias29;
assign weight_bias29= in_buffer_weight29+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias30;
assign weight_bias30= in_buffer_weight30+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias31;
assign weight_bias31= in_buffer_weight31+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias32;
assign weight_bias32= in_buffer_weight32+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias33;
assign weight_bias33= in_buffer_weight33+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias34;
assign weight_bias34= in_buffer_weight34+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias35;
assign weight_bias35= in_buffer_weight35+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias36;
assign weight_bias36= in_buffer_weight36+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias37;
assign weight_bias37= in_buffer_weight37+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias38;
assign weight_bias38= in_buffer_weight38+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias39;
assign weight_bias39= in_buffer_weight39+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias40;
assign weight_bias40= in_buffer_weight40+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias41;
assign weight_bias41= in_buffer_weight41+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias42;
assign weight_bias42= in_buffer_weight42+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias43;
assign weight_bias43= in_buffer_weight43+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias44;
assign weight_bias44= in_buffer_weight44+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias45;
assign weight_bias45= in_buffer_weight45+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias46;
assign weight_bias46= in_buffer_weight46+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias47;
assign weight_bias47= in_buffer_weight47+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias48;
assign weight_bias48= in_buffer_weight48+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias49;
assign weight_bias49= in_buffer_weight49+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias50;
assign weight_bias50= in_buffer_weight50+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias51;
assign weight_bias51= in_buffer_weight51+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias52;
assign weight_bias52= in_buffer_weight52+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias53;
assign weight_bias53= in_buffer_weight53+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias54;
assign weight_bias54= in_buffer_weight54+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias55;
assign weight_bias55= in_buffer_weight55+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias56;
assign weight_bias56= in_buffer_weight56+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias57;
assign weight_bias57= in_buffer_weight57+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias58;
assign weight_bias58= in_buffer_weight58+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias59;
assign weight_bias59= in_buffer_weight59+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias60;
assign weight_bias60= in_buffer_weight60+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias61;
assign weight_bias61= in_buffer_weight61+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias62;
assign weight_bias62= in_buffer_weight62+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias63;
assign weight_bias63= in_buffer_weight63+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias64;
assign weight_bias64= in_buffer_weight64+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias65;
assign weight_bias65= in_buffer_weight65+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias66;
assign weight_bias66= in_buffer_weight66+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias67;
assign weight_bias67= in_buffer_weight67+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias68;
assign weight_bias68= in_buffer_weight68+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias69;
assign weight_bias69= in_buffer_weight69+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias70;
assign weight_bias70= in_buffer_weight70+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias71;
assign weight_bias71= in_buffer_weight71+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias72;
assign weight_bias72= in_buffer_weight72+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias73;
assign weight_bias73= in_buffer_weight73+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias74;
assign weight_bias74= in_buffer_weight74+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias75;
assign weight_bias75= in_buffer_weight75+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias76;
assign weight_bias76= in_buffer_weight76+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias77;
assign weight_bias77= in_buffer_weight77+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias78;
assign weight_bias78= in_buffer_weight78+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias79;
assign weight_bias79= in_buffer_weight79+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias80;
assign weight_bias80= in_buffer_weight80+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias81;
assign weight_bias81= in_buffer_weight81+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias82;
assign weight_bias82= in_buffer_weight82+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias83;
assign weight_bias83= in_buffer_weight83+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias84;
assign weight_bias84= in_buffer_weight84+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias85;
assign weight_bias85= in_buffer_weight85+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias86;
assign weight_bias86= in_buffer_weight86+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias87;
assign weight_bias87= in_buffer_weight87+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias88;
assign weight_bias88= in_buffer_weight88+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias89;
assign weight_bias89= in_buffer_weight89+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias90;
assign weight_bias90= in_buffer_weight90+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias91;
assign weight_bias91= in_buffer_weight91+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias92;
assign weight_bias92= in_buffer_weight92+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias93;
assign weight_bias93= in_buffer_weight93+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias94;
assign weight_bias94= in_buffer_weight94+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias95;
assign weight_bias95= in_buffer_weight95+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias96;
assign weight_bias96= in_buffer_weight96+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias97;
assign weight_bias97= in_buffer_weight97+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias98;
assign weight_bias98= in_buffer_weight98+1;
wire signed    [DATA_WIDTH-1:0]   weight_bias99;
assign weight_bias99= in_buffer_weight99+1;
wire signed    [DATA_WIDTH-1:0]   bias_relu0;
wire signed    [DATA_WIDTH-1:0]   bias_relu1;
wire signed    [DATA_WIDTH-1:0]   bias_relu2;
wire signed    [DATA_WIDTH-1:0]   bias_relu3;
wire signed    [DATA_WIDTH-1:0]   bias_relu4;
wire signed    [DATA_WIDTH-1:0]   bias_relu5;
wire signed    [DATA_WIDTH-1:0]   bias_relu6;
wire signed    [DATA_WIDTH-1:0]   bias_relu7;
wire signed    [DATA_WIDTH-1:0]   bias_relu8;
wire signed    [DATA_WIDTH-1:0]   bias_relu9;
wire signed    [DATA_WIDTH-1:0]   bias_relu10;
wire signed    [DATA_WIDTH-1:0]   bias_relu11;
wire signed    [DATA_WIDTH-1:0]   bias_relu12;
wire signed    [DATA_WIDTH-1:0]   bias_relu13;
wire signed    [DATA_WIDTH-1:0]   bias_relu14;
wire signed    [DATA_WIDTH-1:0]   bias_relu15;
wire signed    [DATA_WIDTH-1:0]   bias_relu16;
wire signed    [DATA_WIDTH-1:0]   bias_relu17;
wire signed    [DATA_WIDTH-1:0]   bias_relu18;
wire signed    [DATA_WIDTH-1:0]   bias_relu19;
wire signed    [DATA_WIDTH-1:0]   bias_relu20;
wire signed    [DATA_WIDTH-1:0]   bias_relu21;
wire signed    [DATA_WIDTH-1:0]   bias_relu22;
wire signed    [DATA_WIDTH-1:0]   bias_relu23;
wire signed    [DATA_WIDTH-1:0]   bias_relu24;
wire signed    [DATA_WIDTH-1:0]   bias_relu25;
wire signed    [DATA_WIDTH-1:0]   bias_relu26;
wire signed    [DATA_WIDTH-1:0]   bias_relu27;
wire signed    [DATA_WIDTH-1:0]   bias_relu28;
wire signed    [DATA_WIDTH-1:0]   bias_relu29;
wire signed    [DATA_WIDTH-1:0]   bias_relu30;
wire signed    [DATA_WIDTH-1:0]   bias_relu31;
wire signed    [DATA_WIDTH-1:0]   bias_relu32;
wire signed    [DATA_WIDTH-1:0]   bias_relu33;
wire signed    [DATA_WIDTH-1:0]   bias_relu34;
wire signed    [DATA_WIDTH-1:0]   bias_relu35;
wire signed    [DATA_WIDTH-1:0]   bias_relu36;
wire signed    [DATA_WIDTH-1:0]   bias_relu37;
wire signed    [DATA_WIDTH-1:0]   bias_relu38;
wire signed    [DATA_WIDTH-1:0]   bias_relu39;
wire signed    [DATA_WIDTH-1:0]   bias_relu40;
wire signed    [DATA_WIDTH-1:0]   bias_relu41;
wire signed    [DATA_WIDTH-1:0]   bias_relu42;
wire signed    [DATA_WIDTH-1:0]   bias_relu43;
wire signed    [DATA_WIDTH-1:0]   bias_relu44;
wire signed    [DATA_WIDTH-1:0]   bias_relu45;
wire signed    [DATA_WIDTH-1:0]   bias_relu46;
wire signed    [DATA_WIDTH-1:0]   bias_relu47;
wire signed    [DATA_WIDTH-1:0]   bias_relu48;
wire signed    [DATA_WIDTH-1:0]   bias_relu49;
wire signed    [DATA_WIDTH-1:0]   bias_relu50;
wire signed    [DATA_WIDTH-1:0]   bias_relu51;
wire signed    [DATA_WIDTH-1:0]   bias_relu52;
wire signed    [DATA_WIDTH-1:0]   bias_relu53;
wire signed    [DATA_WIDTH-1:0]   bias_relu54;
wire signed    [DATA_WIDTH-1:0]   bias_relu55;
wire signed    [DATA_WIDTH-1:0]   bias_relu56;
wire signed    [DATA_WIDTH-1:0]   bias_relu57;
wire signed    [DATA_WIDTH-1:0]   bias_relu58;
wire signed    [DATA_WIDTH-1:0]   bias_relu59;
wire signed    [DATA_WIDTH-1:0]   bias_relu60;
wire signed    [DATA_WIDTH-1:0]   bias_relu61;
wire signed    [DATA_WIDTH-1:0]   bias_relu62;
wire signed    [DATA_WIDTH-1:0]   bias_relu63;
wire signed    [DATA_WIDTH-1:0]   bias_relu64;
wire signed    [DATA_WIDTH-1:0]   bias_relu65;
wire signed    [DATA_WIDTH-1:0]   bias_relu66;
wire signed    [DATA_WIDTH-1:0]   bias_relu67;
wire signed    [DATA_WIDTH-1:0]   bias_relu68;
wire signed    [DATA_WIDTH-1:0]   bias_relu69;
wire signed    [DATA_WIDTH-1:0]   bias_relu70;
wire signed    [DATA_WIDTH-1:0]   bias_relu71;
wire signed    [DATA_WIDTH-1:0]   bias_relu72;
wire signed    [DATA_WIDTH-1:0]   bias_relu73;
wire signed    [DATA_WIDTH-1:0]   bias_relu74;
wire signed    [DATA_WIDTH-1:0]   bias_relu75;
wire signed    [DATA_WIDTH-1:0]   bias_relu76;
wire signed    [DATA_WIDTH-1:0]   bias_relu77;
wire signed    [DATA_WIDTH-1:0]   bias_relu78;
wire signed    [DATA_WIDTH-1:0]   bias_relu79;
wire signed    [DATA_WIDTH-1:0]   bias_relu80;
wire signed    [DATA_WIDTH-1:0]   bias_relu81;
wire signed    [DATA_WIDTH-1:0]   bias_relu82;
wire signed    [DATA_WIDTH-1:0]   bias_relu83;
wire signed    [DATA_WIDTH-1:0]   bias_relu84;
wire signed    [DATA_WIDTH-1:0]   bias_relu85;
wire signed    [DATA_WIDTH-1:0]   bias_relu86;
wire signed    [DATA_WIDTH-1:0]   bias_relu87;
wire signed    [DATA_WIDTH-1:0]   bias_relu88;
wire signed    [DATA_WIDTH-1:0]   bias_relu89;
wire signed    [DATA_WIDTH-1:0]   bias_relu90;
wire signed    [DATA_WIDTH-1:0]   bias_relu91;
wire signed    [DATA_WIDTH-1:0]   bias_relu92;
wire signed    [DATA_WIDTH-1:0]   bias_relu93;
wire signed    [DATA_WIDTH-1:0]   bias_relu94;
wire signed    [DATA_WIDTH-1:0]   bias_relu95;
wire signed    [DATA_WIDTH-1:0]   bias_relu96;
wire signed    [DATA_WIDTH-1:0]   bias_relu97;
wire signed    [DATA_WIDTH-1:0]   bias_relu98;
wire signed    [DATA_WIDTH-1:0]   bias_relu99;
assign bias_relu0=(weight_bias0[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias0;
assign bias_relu1=(weight_bias1[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias1;
assign bias_relu2=(weight_bias2[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias2;
assign bias_relu3=(weight_bias3[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias3;
assign bias_relu4=(weight_bias4[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias4;
assign bias_relu5=(weight_bias5[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias5;
assign bias_relu6=(weight_bias6[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias6;
assign bias_relu7=(weight_bias7[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias7;
assign bias_relu8=(weight_bias8[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias8;
assign bias_relu9=(weight_bias9[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias9;
assign bias_relu10=(weight_bias10[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias10;
assign bias_relu11=(weight_bias11[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias11;
assign bias_relu12=(weight_bias12[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias12;
assign bias_relu13=(weight_bias13[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias13;
assign bias_relu14=(weight_bias14[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias14;
assign bias_relu15=(weight_bias15[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias15;
assign bias_relu16=(weight_bias16[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias16;
assign bias_relu17=(weight_bias17[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias17;
assign bias_relu18=(weight_bias18[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias18;
assign bias_relu19=(weight_bias19[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias19;
assign bias_relu20=(weight_bias20[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias20;
assign bias_relu21=(weight_bias21[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias21;
assign bias_relu22=(weight_bias22[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias22;
assign bias_relu23=(weight_bias23[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias23;
assign bias_relu24=(weight_bias24[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias24;
assign bias_relu25=(weight_bias25[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias25;
assign bias_relu26=(weight_bias26[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias26;
assign bias_relu27=(weight_bias27[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias27;
assign bias_relu28=(weight_bias28[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias28;
assign bias_relu29=(weight_bias29[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias29;
assign bias_relu30=(weight_bias30[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias30;
assign bias_relu31=(weight_bias31[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias31;
assign bias_relu32=(weight_bias32[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias32;
assign bias_relu33=(weight_bias33[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias33;
assign bias_relu34=(weight_bias34[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias34;
assign bias_relu35=(weight_bias35[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias35;
assign bias_relu36=(weight_bias36[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias36;
assign bias_relu37=(weight_bias37[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias37;
assign bias_relu38=(weight_bias38[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias38;
assign bias_relu39=(weight_bias39[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias39;
assign bias_relu40=(weight_bias40[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias40;
assign bias_relu41=(weight_bias41[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias41;
assign bias_relu42=(weight_bias42[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias42;
assign bias_relu43=(weight_bias43[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias43;
assign bias_relu44=(weight_bias44[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias44;
assign bias_relu45=(weight_bias45[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias45;
assign bias_relu46=(weight_bias46[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias46;
assign bias_relu47=(weight_bias47[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias47;
assign bias_relu48=(weight_bias48[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias48;
assign bias_relu49=(weight_bias49[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias49;
assign bias_relu50=(weight_bias50[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias50;
assign bias_relu51=(weight_bias51[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias51;
assign bias_relu52=(weight_bias52[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias52;
assign bias_relu53=(weight_bias53[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias53;
assign bias_relu54=(weight_bias54[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias54;
assign bias_relu55=(weight_bias55[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias55;
assign bias_relu56=(weight_bias56[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias56;
assign bias_relu57=(weight_bias57[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias57;
assign bias_relu58=(weight_bias58[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias58;
assign bias_relu59=(weight_bias59[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias59;
assign bias_relu60=(weight_bias60[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias60;
assign bias_relu61=(weight_bias61[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias61;
assign bias_relu62=(weight_bias62[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias62;
assign bias_relu63=(weight_bias63[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias63;
assign bias_relu64=(weight_bias64[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias64;
assign bias_relu65=(weight_bias65[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias65;
assign bias_relu66=(weight_bias66[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias66;
assign bias_relu67=(weight_bias67[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias67;
assign bias_relu68=(weight_bias68[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias68;
assign bias_relu69=(weight_bias69[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias69;
assign bias_relu70=(weight_bias70[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias70;
assign bias_relu71=(weight_bias71[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias71;
assign bias_relu72=(weight_bias72[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias72;
assign bias_relu73=(weight_bias73[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias73;
assign bias_relu74=(weight_bias74[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias74;
assign bias_relu75=(weight_bias75[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias75;
assign bias_relu76=(weight_bias76[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias76;
assign bias_relu77=(weight_bias77[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias77;
assign bias_relu78=(weight_bias78[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias78;
assign bias_relu79=(weight_bias79[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias79;
assign bias_relu80=(weight_bias80[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias80;
assign bias_relu81=(weight_bias81[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias81;
assign bias_relu82=(weight_bias82[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias82;
assign bias_relu83=(weight_bias83[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias83;
assign bias_relu84=(weight_bias84[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias84;
assign bias_relu85=(weight_bias85[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias85;
assign bias_relu86=(weight_bias86[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias86;
assign bias_relu87=(weight_bias87[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias87;
assign bias_relu88=(weight_bias88[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias88;
assign bias_relu89=(weight_bias89[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias89;
assign bias_relu90=(weight_bias90[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias90;
assign bias_relu91=(weight_bias91[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias91;
assign bias_relu92=(weight_bias92[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias92;
assign bias_relu93=(weight_bias93[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias93;
assign bias_relu94=(weight_bias94[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias94;
assign bias_relu95=(weight_bias95[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias95;
assign bias_relu96=(weight_bias96[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias96;
assign bias_relu97=(weight_bias97[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias97;
assign bias_relu98=(weight_bias98[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias98;
assign bias_relu99=(weight_bias99[DATA_WIDTH-1]==1'b1)   ?   {DATA_WIDTH{1'b0}}:weight_bias99;
assign layer_out={
bias_relu99,bias_relu98,bias_relu97,bias_relu96,bias_relu95,bias_relu94,bias_relu93,bias_relu92,bias_relu91,bias_relu90,bias_relu89,bias_relu88,bias_relu87,bias_relu86,bias_relu85,bias_relu84,bias_relu83,bias_relu82,bias_relu81,bias_relu80,bias_relu79,bias_relu78,bias_relu77,bias_relu76,bias_relu75,bias_relu74,bias_relu73,bias_relu72,bias_relu71,bias_relu70,bias_relu69,bias_relu68,bias_relu67,bias_relu66,bias_relu65,bias_relu64,bias_relu63,bias_relu62,bias_relu61,bias_relu60,bias_relu59,bias_relu58,bias_relu57,bias_relu56,bias_relu55,bias_relu54,bias_relu53,bias_relu52,bias_relu51,bias_relu50,bias_relu49,bias_relu48,bias_relu47,bias_relu46,bias_relu45,bias_relu44,bias_relu43,bias_relu42,bias_relu41,bias_relu40,bias_relu39,bias_relu38,bias_relu37,bias_relu36,bias_relu35,bias_relu34,bias_relu33,bias_relu32,bias_relu31,bias_relu30,bias_relu29,bias_relu28,bias_relu27,bias_relu26,bias_relu25,bias_relu24,bias_relu23,bias_relu22,bias_relu21,bias_relu20,bias_relu19,bias_relu18,bias_relu17,bias_relu16,bias_relu15,bias_relu14,bias_relu13,bias_relu12,bias_relu11,bias_relu10,bias_relu9,bias_relu8,bias_relu7,bias_relu6,bias_relu5,bias_relu4,bias_relu3,bias_relu2,bias_relu1,bias_relu0};
always@(posedge clk)
    begin
        if(rst)
            begin
                ready<=1'b0;
            end
        else
            begin
                ready<=valid;
            end
    end
endmodule